`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:       James Swineson
// 
// Create Date:    14:47:27 12/30/2017 
// Design Name:    ButtonDejitter
// Module Name:    ButtonDejitter.v
// Project Name:   ButtonDejitter
// Target Devices: XC6LX16
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

// Generated by the following python code:
//   for i in range(1, 32): print("(x <= {})?{}:\\".format(2**i, i))
// we end at 4294967295 since default int is 32 bit.
// use WIDTH'dxxxx if larger int is needed.
// the last -1 is used to indicater no LUT value error.
`define CLOG2(x) \
(x <= 2)?1:\
(x <= 4)?2:\
(x <= 8)?3:\
(x <= 16)?4:\
(x <= 32)?5:\
(x <= 64)?6:\
(x <= 128)?7:\
(x <= 256)?8:\
(x <= 512)?9:\
(x <= 1024)?10:\
(x <= 2048)?11:\
(x <= 4096)?12:\
(x <= 8192)?13:\
(x <= 16384)?14:\
(x <= 32768)?15:\
(x <= 65536)?16:\
(x <= 131072)?17:\
(x <= 262144)?18:\
(x <= 524288)?19:\
(x <= 1048576)?20:\
(x <= 2097152)?21:\
(x <= 4194304)?22:\
(x <= 8388608)?23:\
(x <= 16777216)?24:\
(x <= 33554432)?25:\
(x <= 67108864)?26:\
(x <= 134217728)?27:\
(x <= 268435456)?28:\
(x <= 536870912)?29:\
(x <= 1073741824)?30:\
(x <= 2147483648)?31:\
(x <= 4294967295)?32:\
	-1

module ButtonDejitter #(
		parameter COUNT_TO = 5000000,
		parameter DATA_WIDTH = `CLOG2(COUNT_TO) + 1
	)(
    input BTN_IN,
    input CLK,
    output BTN_OUT
    );

reg DEJITTERED = 0;
reg [DATA_WIDTH:0] count = 0;

assign BTN_OUT = DEJITTERED;

always @(posedge CLK) begin
	if (BTN_IN != DEJITTERED) count = count + 1;
	else count = 0;
	
	if (count == COUNT_TO) begin
		DEJITTERED = BTN_IN;
		count = 0;
	end
end

endmodule
